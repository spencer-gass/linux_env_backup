// CONFIDENTIAL
// Copyright (c) 2024 Kepler Communications Inc.

`timescale 1ns/1ps
`include "../util/util_check_elab.svh"
`default_nettype none

/**
 * Egress subsystem for P4 router
 *  Input wide AXIS bus from VNP4
 *  axis_demux_wrapper to split out to egress port buffers
 *  axis_adapt to width convert
 *  output to physical ports
**/
module p4_router_egress
    import P4_ROUTER_PKG::*;
 #(
    parameter int                               NUM_8B_EGR_PHYS_PORTS  = 0,
    parameter int                               NUM_16B_EGR_PHYS_PORTS = 0,
    parameter int                               NUM_32B_EGR_PHYS_PORTS = 0,
    parameter int                               NUM_64B_EGR_PHYS_PORTS = 0,
    parameter int                               MTU_BYTES              = 1500,
    parameter int                               NUM_EGR_PHYS_PORTS     = NUM_64B_EGR_PHYS_PORTS
                                                                       + NUM_32B_EGR_PHYS_PORTS
                                                                       + NUM_16B_EGR_PHYS_PORTS
                                                                       + NUM_8B_EGR_PHYS_PORTS,

    parameter bit                               EGR_BUS_DEBUG_ILA      = 1'b0,
    parameter bit [NUM_8B_EGR_PHYS_PORTS-1:0]   EGR_8B_PORT_DEBUG_ILA  = '0,
    parameter bit [NUM_16B_EGR_PHYS_PORTS-1:0]  EGR_16B_PORT_DEBUG_ILA = '0,
    parameter bit [NUM_32B_EGR_PHYS_PORTS-1:0]  EGR_32B_PORT_DEBUG_ILA = '0,
    parameter bit [NUM_64B_EGR_PHYS_PORTS-1:0]  EGR_64B_PORT_DEBUG_ILA = '0
)(
    AXIS_int.Slave                            egr_bus,
    output var logic [NUM_EGR_PHYS_PORTS-1:0] egr_buf_ready,

    AXIS_int.Master                           egr_8b_phys_ports  [NUM_8B_EGR_PHYS_PORTS-1:0],  // Can't group interfaces with different parameters into an array. One array per data width supported.
    AXIS_int.Master                           egr_16b_phys_ports [NUM_16B_EGR_PHYS_PORTS-1:0],
    AXIS_int.Master                           egr_32b_phys_ports [NUM_32B_EGR_PHYS_PORTS-1:0],
    AXIS_int.Master                           egr_64b_phys_ports [NUM_64B_EGR_PHYS_PORTS-1:0],

    input  var logic [NUM_EGR_PHYS_PORTS-1:0] egr_phys_ports_enable,
    input  var logic [NUM_EGR_PHYS_PORTS-1:0] egr_cnts_clear,
    output var logic [EGR_COUNTERS_WIDTH-1:0] egr_cnts [NUM_EGR_PHYS_PORTS-1:0] [6:0],
    output var logic [NUM_EGR_PHYS_PORTS-1:0] egr_ports_conneted,
    output var logic [NUM_EGR_PHYS_PORTS-1:0] egr_buf_full_drop
);


    ////////////////////////////////////////////////////////////////////////////////////////////////
    // SECTION: Localparams


    localparam int NUM_EGR_PHYS_PORTS_PER_ARRAY [NUM_EGR_AXIS_ARRAYS-1:0] = {NUM_64B_EGR_PHYS_PORTS,
                                                                             NUM_32B_EGR_PHYS_PORTS,
                                                                             NUM_16B_EGR_PHYS_PORTS,
                                                                             NUM_8B_EGR_PHYS_PORTS
                                                                          };

    localparam int MAX_NUM_PORTS_PER_ARRAY = get_max_num_ports_per_array(NUM_EGR_PHYS_PORTS_PER_ARRAY);

    typedef int egr_port_index_map_t [NUM_EGR_AXIS_ARRAYS-1:0] [MAX_NUM_PORTS_PER_ARRAY-1:0];

    function automatic egr_port_index_map_t create_egr_port_index_map();
        begin
            automatic egr_port_index_map_t map = '{default: '{default: -1}};
            automatic int cnt = 0;
            for(int i=0; i<NUM_EGR_AXIS_ARRAYS; i++) begin
                for(int j=0; j<NUM_EGR_PHYS_PORTS_PER_ARRAY[i]; j++) begin
                    map[i][j] = cnt;
                    cnt++;
                end
            end
            return map;
        end
    endfunction

    localparam NUM_EGR_PHYS_PORTS_LOG = $clog2(NUM_EGR_PHYS_PORTS);

    localparam egr_port_index_map_t EGR_PORT_INDEX_MAP = create_egr_port_index_map();


    ////////////////////////////////////////////////////////////////////////////////////////////////
    // SECTION: Elaboration Checks


    `ELAB_CHECK_GE(egr_bus.DATA_BYTES, 8) // wide output bus needs to be at least as wide as the widest input bus
    `ELAB_CHECK_GT(NUM_EGR_PHYS_PORTS, 0);
    `ELAB_CHECK_EQUAL(NUM_EGR_PHYS_PORTS, NUM_64B_EGR_PHYS_PORTS
                                        + NUM_32B_EGR_PHYS_PORTS
                                        + NUM_16B_EGR_PHYS_PORTS
                                        + NUM_8B_EGR_PHYS_PORTS);


    ////////////////////////////////////////////////////////////////////////////////////////////////
    // SECTION: Signal Declarations


    AXIS_int #(
        .DATA_BYTES ( egr_bus.DATA_BYTES  )
    ) egr_phys_ports_demuxed [NUM_EGR_PHYS_PORTS-1:0] (
        .clk     ( egr_bus.clk     ),
        .sresetn ( egr_bus.sresetn )
    );

    queue_system_metadata_t queue_system_metadata;
    logic [NUM_EGR_PHYS_PORTS_LOG-1:0] egr_port_sel;


    ////////////////////////////////////////////////////////////////////////////////////////////////
    // SECTION: Egress Demux


    assign queue_system_metadata    = egr_bus.tuser;
    assign egr_port_sel             = queue_system_metadata.egress_port[NUM_EGR_PHYS_PORTS_LOG-1:0];
    assign egr_bus.tready           = 1'b1;

    generate
        for (genvar port=0; port<NUM_EGR_PHYS_PORTS; port++) begin : egress_demux
            assign egr_buf_ready[port] = egr_phys_ports_demuxed[port].tready;
            always_ff @(posedge egr_bus.clk) begin
                egr_phys_ports_demuxed[port].tvalid <= (egr_bus.tvalid && egr_port_sel === port && egr_bus.sresetn) ? 1'b1 : 1'b0;
                egr_phys_ports_demuxed[port].tdata  <= egr_bus.tdata;
                egr_phys_ports_demuxed[port].tstrb  <= egr_bus.tstrb;
                egr_phys_ports_demuxed[port].tkeep  <= egr_bus.tkeep;
                egr_phys_ports_demuxed[port].tlast  <= egr_bus.tlast;
                egr_phys_ports_demuxed[port].tid    <= egr_bus.tid;
                egr_phys_ports_demuxed[port].tdest  <= egr_bus.tdest;
                egr_phys_ports_demuxed[port].tuser  <= 1'b0;
            end
        end
    endgenerate



    ////////////////////////////////////////////////////////////////////////////////////////////////
    // SECTION: Per-Physical-Port Logic


    // For each egress physical port, convert data bus width to physical port width

    `define DEF_EGR_PORT_ADAPT(WIDTH, BYTES)                                                                                    \
        p4_router_egress_port_array_adapt #(                                                                                    \
            .NUM_EGR_PHYS_PORTS         ( NUM_``WIDTH``B_EGR_PHYS_PORTS ),                                                      \
            .EGR_BUS_DATA_BYTES         ( egr_bus.DATA_BYTES            ),                                                      \
            .PHYS_PORT_DATA_BYTES       ( BYTES                         ),                                                      \
            .MTU_BYTES                  ( MTU_BYTES                     ),                                                      \
            .EGR_COUNTERS_WIDTH         ( EGR_COUNTERS_WIDTH            )                                                       \
        ) egress_port_array_adapt_``WIDTH``b (                                                                                  \
            .egr_phys_ports_demuxed     ( egr_phys_ports_demuxed[INDEX_``WIDTH``B_START +: NUM_``WIDTH``B_EGR_PHYS_PORTS]   ),  \
            .egr_phys_ports             ( egr_``WIDTH``b_phys_ports                                                         ),  \
            .egr_phys_ports_enable      ( egr_phys_ports_enable [INDEX_``WIDTH``B_START +: NUM_``WIDTH``B_EGR_PHYS_PORTS]   ),  \
            .egr_cnts_clear             ( egr_cnts_clear        [INDEX_``WIDTH``B_START +: NUM_``WIDTH``B_EGR_PHYS_PORTS]   ),  \
            .egr_cnts                   ( egr_cnts              [INDEX_``WIDTH``B_START +: NUM_``WIDTH``B_EGR_PHYS_PORTS]   ),  \
            .egr_ports_connected        ( egr_ports_conneted    [INDEX_``WIDTH``B_START +: NUM_``WIDTH``B_EGR_PHYS_PORTS]   ),  \
            .egr_buf_full_drop          ( egr_buf_full_drop     [INDEX_``WIDTH``B_START +: NUM_``WIDTH``B_EGR_PHYS_PORTS]   )   \
        );
    generate
        if (NUM_8B_EGR_PHYS_PORTS) begin : adapt_8b
            `DEF_EGR_PORT_ADAPT(8, 1);
        end

        if (NUM_16B_EGR_PHYS_PORTS) begin : adapt_16b
            `DEF_EGR_PORT_ADAPT(16, 2);
        end

        if (NUM_32B_EGR_PHYS_PORTS) begin : adapt_32b
            `DEF_EGR_PORT_ADAPT(32, 4);
        end

        if (NUM_64B_EGR_PHYS_PORTS) begin : adapt_64b
            `DEF_EGR_PORT_ADAPT(64, 8);
        end
    endgenerate

    `ifndef MODEL_TECH
        /* svlint off style_keyword_end */
        `define DEF_EGR_PORT_ILA(WIDTH)                                     \
            logic [31:0] dbg_cntr;                                          \
            always_ff @(posedge egr_``WIDTH``b_phys_ports[port].clk) begin  \
                if (!egr_``WIDTH``b_phys_ports[port].sresetn) begin         \
                    dbg_cntr <= '0;                                         \
                end else begin                                              \
                    dbg_cntr <= dbg_cntr + 1'b1;                            \
                end                                                         \
            end                                                             \
                                                                            \
            ila_debug egr_``WIDTH``b_port_ila (                             \
                .clk    ( egr_``WIDTH``b_phys_ports[port].clk       ),      \
                .probe0 ( egr_``WIDTH``b_phys_ports[port].sresetn   ),      \
                .probe1 ( egr_``WIDTH``b_phys_ports[port].tready    ),      \
                .probe2 ( egr_``WIDTH``b_phys_ports[port].tvalid    ),      \
                .probe3 ( egr_``WIDTH``b_phys_ports[port].tdata     ),      \
                .probe4 ( egr_``WIDTH``b_phys_ports[port].tkeep     ),      \
                .probe5 ( egr_``WIDTH``b_phys_ports[port].tlast     ),      \
                .probe6 ( dbg_cntr                                  ),      \
                .probe7 ( '0                                        ),      \
                .probe8 ( '0                                        ),      \
                .probe9 ( '0                                        ),      \
                .probe10( '0                                        ),      \
                .probe11( '0                                        ),      \
                .probe12( '0                                        ),      \
                .probe13( '0                                        ),      \
                .probe14( '0                                        ),      \
                .probe15( '0                                        )       \
            );

        generate
                if (EGR_BUS_DEBUG_ILA) begin : gen_ila
                    logic [31:0] dbg_cntr;
                    always_ff @(posedge egr_bus.clk) begin
                        if (!egr_bus.sresetn) begin
                            dbg_cntr <= '0;
                        end else begin
                            dbg_cntr <= dbg_cntr + 1'b1;
                        end
                    end

                    ila_debug egr_bus_ila (
                        .clk    ( egr_bus.clk       ),
                        .probe0 ( egr_bus.sresetn   ),
                        .probe1 ( egr_bus.tready    ),
                        .probe2 ( egr_bus.tvalid    ),
                        .probe3 ( egr_bus.tkeep     ),
                        .probe4 ( egr_bus.tlast     ),
                        .probe5 ( egr_bus.tuser     ),
                        .probe6 ( dbg_cntr          ),
                        .probe7 ( '0                ),
                        .probe8 ( '0                ),
                        .probe9 ( '0                ),
                        .probe10( '0                ),
                        .probe11( '0                ),
                        .probe12( '0                ),
                        .probe13( '0                ),
                        .probe14( '0                ),
                        .probe15( '0                )
                    );
                end


            for (genvar port=0; port<NUM_8B_EGR_PHYS_PORTS; port++) begin : ila_8b
                if (EGR_8B_PORT_DEBUG_ILA[port]) begin : gen_ila
                    `DEF_EGR_PORT_ILA(8);
                end
            end

            for (genvar port=0; port<NUM_16B_EGR_PHYS_PORTS; port++) begin : ila_16b
                if (EGR_16B_PORT_DEBUG_ILA[port]) begin : gen_ila
                    `DEF_EGR_PORT_ILA(16);
                end
            end

            for (genvar port=0; port<NUM_32B_EGR_PHYS_PORTS; port++) begin : ila_32b
                if (EGR_32B_PORT_DEBUG_ILA[port]) begin : gen_ila
                    `DEF_EGR_PORT_ILA(32);
                end
            end

            for (genvar port=0; port<NUM_64B_EGR_PHYS_PORTS; port++) begin : ila_64b
                if (EGR_64B_PORT_DEBUG_ILA[port]) begin : gen_ila
                    `DEF_EGR_PORT_ILA(64);
                end
            end
        endgenerate
    `endif
    /* svlint on style_keyword_end */

endmodule

`default_nettype wire
