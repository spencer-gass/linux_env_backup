// CONFIDENTIAL
// Copyright (c) 2024 Kepler Communications Inc.

/**
 * IPv4 Check Sum Test Bench Package
**/

`default_nettype none

package ipv4_checksum_tb_pkg;

    ////////////////////////////////////////////////////////////////////////////////////////////////
    // SECTION: Imports

    ////////////////////////////////////////////////////////////////////////////////////////////////
    // SECTION: Localparams


    ////////////////////////////////////////////////////////////////////////////////////////////////
    // SECTION: Type Definitions

    ////////////////////////////////////////////////////////////////////////////////////////////////
    // SECTION: Functions


endpackage