// CONFIDENTIAL
// Copyright (c) 2024 Kepler Communications Inc.

/**
 * Encapsulate packet gens into a module so that there can be one perameterized module instantiatoin per
 * axis array ranther than four instances of nearly identical logic.
 */

`include "../../rtl/util/util_check_elab.svh"
`default_nettype none
`timescale 1ns/1ps

module axis_array_packet_generator
#(
    parameter NUM_PORTS = 0,
    parameter MTU_BYTES = 1500

) (
    AXIS_int.Master axis_packet_out [NUM_PORTS-1:0],

    output var logic [NUM_PORTS-1:0]                        busy,
    input  var logic [NUM_PORTS-1:0]                        send_packet_req,
    input  var int                                          packet_byte_length  [NUM_PORTS-1:0],
    input  var logic [axis_packet_out[0].USER_WIDTH-1:0]    packet_user         [NUM_PORTS-1:0],
    input  var logic [MTU_BYTES*8-1:0]                      packet_data         [NUM_PORTS-1:0]
);

    `ELAB_CHECK_GT(NUM_PORTS, 0);

    generate
        for (genvar port=0; port < NUM_PORTS; port++) begin
            axis_packet_generator #(
                .MTU_BYTES (MTU_BYTES)
            ) packet_generator (
                .axis_packet_out     ( axis_packet_out[port]    ),
                .busy                ( busy[port]               ),
                .send_packet_req     ( send_packet_req[port]    ),
                .packet_byte_length  ( packet_byte_length[port] ),
                .packet_user         ( packet_user[port]        ),
                .packet_data         ( packet_data[port]        )
            );
        end
    endgenerate

endmodule
