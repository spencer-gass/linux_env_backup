// CONFIDENTIAL
// Copyright (c) 2024 Kepler Communications Inc.

`include "vunit_defines.svh"
`include "../../rtl/util/util_check_elab.svh"
`include "../../rtl/util/util_make_monitors.svh"
`default_nettype none
`timescale 1ns/1ps

/**
 * Test bench for p4_router_egress.
 */
module p4_router_egress_tb ();


    ////////////////////////////////////////////////////////////////////////////////////////////////
    // SECTION: Parameter definition


    parameter int NUM_8B_PORTS          = 3;    // Number of 8-bit  physical ports to the DUT
    parameter int NUM_16B_PORTS         = 0;    // Number of 16-bit physical ports to the DUT
    parameter int NUM_32B_PORTS         = 3;    // Number of 32-bit physical ports to the DUT
    parameter int NUM_64B_PORTS         = 0;    // Number of 640bit physical ports to the DUT
    parameter int EGR_AXIS_DATA_BYTES   = 8;    // Width of axis bus toward VNP4
    parameter int MTU_BYTES             = 1500; // MTU for the router
    parameter int PACKET_MAX_BLEN       = 1000; // Maximum packet size in BYTES
    parameter int PACKET_MIN_BLEN       = 64;   // Minimum packet size in BYTES
    parameter int NUM_PACKETS_TO_SEND   = 100;


    ////////////////////////////////////////////////////////////////////////////////////////////////
    // SECTION: Import


    import P4_ROUTER_PKG::*;
    import P4_ROUTER_TB_PKG::*;
    import UTIL_INTS::U_INT_CEIL_DIV;


    ////////////////////////////////////////////////////////////////////////////////////////////////
    // SECTION: Constants


    localparam int PAYLOAD_TYPE = RAND;

    localparam int NUM_EGR_PHYS_PORTS_PER_ARRAY [NUM_EGR_AXIS_ARRAYS-1:0] = {NUM_64B_PORTS,
                                                                             NUM_32B_PORTS,
                                                                             NUM_16B_PORTS,
                                                                             NUM_8B_PORTS
                                                                          };

    localparam int NUM_PORTS      = NUM_8B_PORTS + NUM_16B_PORTS + NUM_32B_PORTS + NUM_64B_PORTS;
    localparam int NUM_PORTS_LOG  = $clog2(NUM_PORTS);

    localparam port_index_map_t EGR_PORT_INDEX_MAP = create_port_index_map(NUM_EGR_PHYS_PORTS_PER_ARRAY);

    localparam int EGR_8B_START  = EGR_PORT_INDEX_MAP[INDEX_8B][0];
    localparam int EGR_16B_START = EGR_PORT_INDEX_MAP[INDEX_16B][0];
    localparam int EGR_32B_START = EGR_PORT_INDEX_MAP[INDEX_32B][0];
    localparam int EGR_64B_START = EGR_PORT_INDEX_MAP[INDEX_64B][0];

    localparam int MAX_PKT_EGR_WLEN = U_INT_CEIL_DIV(PACKET_MAX_BLEN, EGR_AXIS_DATA_BYTES);
    localparam int MAX_PKT_WLEN_8B  = PACKET_MAX_BLEN/BYTES_PER_8BIT_WORD;

    localparam int MTU_BYTES_LOG            = $clog2(MTU_BYTES);
    localparam int NUM_PACKETS_TO_SEND_LOG  = $clog2(NUM_PACKETS_TO_SEND);


    ////////////////////////////////////////////////////////////////////////////////////////////////
    // SECTION: Signal Declarations


    bit   [NUM_PORTS-1:0]           egr_buf_ready;
    bit   [NUM_PORTS-1:0]           egr_phys_ports_enable;
    bit   [NUM_PORTS-1:0]           egr_cnts_clear;
    logic [EGR_COUNTERS_WIDTH-1:0]  egr_cnts [NUM_PORTS-1:0] [6:0];
    bit   [NUM_PORTS-1:0]           egr_ports_conneted;

    int                             send_packet_byte_length;
    queue_system_metadata_t         send_packet_user;

    logic [0:MTU_BYTES*8-1]         send_packet_data;
    bit                             send_packet_req;
    bit                             send_packet_req_d;
    bit   [NUM_PORTS-1:0]           send_packet_busy;

    int   expected_count;
    int   received_count_array [NUM_PORTS-1:0];
    int   received_count;
    bit   packet_received;

    bit   [NUM_PORTS-1:0] egr_phys_ports_tlast;
    bit   [NUM_PORTS-1:0] egr_phys_ports_tvalid;

    bit   [EGR_COUNTERS_WIDTH-1:0] expected_egr_cnts [NUM_PORTS-1:0] [6:0];

    bit   [NUM_PORTS-1:0]  egr_buf_full_drop;
    bit   [NUM_PORTS-1:0]  egr_buf_full_drop_sticky;
    bit                    egr_buf_full_drop_clear;

    bit   verify_sequence;
    int   seq_cnt;

    logic [0:MTU_BYTES*8-1]             tx_snoop_data_buf   [NUM_PORTS-1:0] [NUM_PACKETS_TO_SEND-1:0];
    logic [MTU_BYTES_LOG-1:0]           tx_snoop_blen_buf   [NUM_PORTS-1:0] [NUM_PACKETS_TO_SEND-1:0];
    logic [NUM_PACKETS_TO_SEND_LOG:0]   tx_snoop_wr_ptr     [NUM_PORTS-1:0];

    logic [0:MTU_BYTES*8-1]     send_data_buf        [NUM_PORTS-1:0];
    int                         send_byte_length_buf [NUM_PORTS-1:0];
    queue_system_metadata_t     send_user_buf        [NUM_PORTS-1:0];
    int                         send_egr_port;
    int                         egr_port_rr;

    bit   [EGR_AXIS_DATA_BYTES-1:0] tkeep_comb;

    bit   [NUM_8B_PORTS-1:0]  egr_8b_async_fifo_overflow  = '0;
    bit   [NUM_16B_PORTS-1:0] egr_16b_async_fifo_overflow = '0;
    bit   [NUM_32B_PORTS-1:0] egr_32b_async_fifo_overflow = '0;
    bit   [NUM_64B_PORTS-1:0] egr_64b_async_fifo_overflow = '0;

    logic [DQ_LATENCY-1:0] dq_in_flight [NUM_PORTS-1:0];


    ////////////////////////////////////////////////////////////////////////////////////////////////
    // SECTION: AXIS Declarations


    AXIS_int #(
        .DATA_BYTES ( EGR_AXIS_DATA_BYTES           ),
        .USER_WIDTH ( VNP4_WRAPPER_METADATA_WIDTH   )
    ) egr_bus (
        .clk     (core_clk_ifc.clk                                      ),
        .sresetn (core_sreset_ifc.reset != core_sreset_ifc.ACTIVE_HIGH  )
    );

    AXIS_int #(
        .DATA_BYTES ( BYTES_PER_8BIT_WORD )
    ) egr_8b_phys_ports [NUM_8B_PORTS-1:0] (
        .clk     (core_clk_ifc.clk                                      ),
        .sresetn (core_sreset_ifc.reset != core_sreset_ifc.ACTIVE_HIGH  )
    );

    AXIS_int #(
        .DATA_BYTES ( BYTES_PER_16BIT_WORD )
    ) egr_16b_phys_ports [NUM_16B_PORTS-1:0] (
        .clk     (core_clk_ifc.clk                                      ),
        .sresetn (core_sreset_ifc.reset != core_sreset_ifc.ACTIVE_HIGH  )
    );

    AXIS_int #(
        .DATA_BYTES ( BYTES_PER_32BIT_WORD )
    ) egr_32b_phys_ports [NUM_32B_PORTS-1:0] (
        .clk     (core_clk_ifc.clk                                      ),
        .sresetn (core_sreset_ifc.reset != core_sreset_ifc.ACTIVE_HIGH  )
    );

    AXIS_int #(
        .DATA_BYTES ( BYTES_PER_64BIT_WORD )
    ) egr_64b_phys_ports [NUM_64B_PORTS-1:0] (
        .clk     (core_clk_ifc.clk                                      ),
        .sresetn (core_sreset_ifc.reset != core_sreset_ifc.ACTIVE_HIGH  )
    );

    AXIS_int #(
        .DATA_BYTES ( BYTES_PER_8BIT_WORD )
    ) egr_8b_phys_ports_cdc [NUM_8B_PORTS-1:0] (
        .clk     (egr_port_clk_ifc.clk                                         ),
        .sresetn (egr_port_sreset_ifc.reset != egr_port_sreset_ifc.ACTIVE_HIGH )
    );

    AXIS_int #(
        .DATA_BYTES ( BYTES_PER_16BIT_WORD )
    ) egr_16b_phys_ports_cdc [NUM_16B_PORTS-1:0] (
        .clk     (egr_port_clk_ifc.clk                                         ),
        .sresetn (egr_port_sreset_ifc.reset != egr_port_sreset_ifc.ACTIVE_HIGH )
    );

    AXIS_int #(
        .DATA_BYTES ( BYTES_PER_32BIT_WORD )
    ) egr_32b_phys_ports_cdc [NUM_32B_PORTS-1:0] (
        .clk     (egr_port_clk_ifc.clk                                         ),
        .sresetn (egr_port_sreset_ifc.reset != egr_port_sreset_ifc.ACTIVE_HIGH )
    );

    AXIS_int #(
        .DATA_BYTES ( BYTES_PER_64BIT_WORD )
    ) egr_64b_phys_ports_cdc [NUM_64B_PORTS-1:0] (
        .clk     (egr_port_clk_ifc.clk                                         ),
        .sresetn (egr_port_sreset_ifc.reset != egr_port_sreset_ifc.ACTIVE_HIGH )
    );

    Clock_int #(
        .CLOCK_GROUP_ID   ( 0 ),
        .SOURCE_FREQUENCY ( 0 )
    ) egr_port_clk_ifc ();

    Reset_int #(
        .CLOCK_GROUP_ID ( 0 )
    ) egr_port_sreset_ifc ();

    Clock_int #(
        .CLOCK_GROUP_ID   ( 0 ),
        .SOURCE_FREQUENCY ( 0 )
    ) core_clk_ifc ();

    Reset_int #(
        .CLOCK_GROUP_ID ( 0 )
    ) core_sreset_ifc ();


    ////////////////////////////////////////////////////////////////////////////////////////////////
    // SECTION: Logic Implemenatation


    // Simulation Clocks
    always #(PHYS_PORT_CLK_PERIOD/2) egr_port_clk_ifc.clk <= ~egr_port_clk_ifc.clk;
    always #(CORE_CLK_PERIOD/2)      core_clk_ifc.clk     <= ~core_clk_ifc.clk;


    ////////////////////////////////////////////////////////////////////////////////////////////////
    // SUB-SECTION: Packet Generator


    assign send_egr_port = send_packet_user.egress_port[NUM_PORTS_LOG-1:0];

    always_comb begin
        for (int port=0; port<NUM_PORTS; port++) begin
            send_packet_busy[port] = (send_byte_length_buf[port] === 0) ? 1'b0 : 1'b1;
        end
    end

    always_comb begin
        tkeep_comb = '0;
        for (int b=0; b<EGR_AXIS_DATA_BYTES; b++) begin
            if (send_byte_length_buf[egr_port_rr] % EGR_AXIS_DATA_BYTES == 0) begin
                tkeep_comb[b] = 1'b1;
            end else if (b < send_byte_length_buf[egr_port_rr] % EGR_AXIS_DATA_BYTES) begin
                tkeep_comb[b] = 1'b1;
            end
        end
    end

    always_ff @(posedge core_clk_ifc.clk) begin
        if (core_sreset_ifc.reset == core_sreset_ifc.ACTIVE_HIGH) begin
            send_data_buf        <= '{default: '0};
            send_byte_length_buf <= '{default: 0};
            send_user_buf        <= '{default: '0};
            egr_port_rr          <= 0;
            dq_in_flight         <= '{default: '0};
        end else begin
            if (send_packet_req && !send_packet_req_d && !send_packet_busy[send_egr_port]) begin
                send_data_buf[send_egr_port]        <= send_packet_data;
                send_byte_length_buf[send_egr_port] <= send_packet_byte_length;
                send_user_buf[send_egr_port]        <= send_packet_user;
            end

            if (egr_port_rr == NUM_PORTS-1) begin
                egr_port_rr <= 0;
            end else begin
                egr_port_rr <= egr_port_rr + 1;
            end

            for (int port=0; port<NUM_PORTS; port++) begin
                dq_in_flight[port] <= {dq_in_flight[port][DQ_LATENCY-2:0], 1'b0};
            end

            egr_bus.tlast  <= 1'b0;
            egr_bus.tkeep  <= '1;
            egr_bus.tvalid <= 1'b0;
            if (egr_buf_ready[egr_port_rr] && send_packet_busy[egr_port_rr] && ~|dq_in_flight[egr_port_rr]) begin
                egr_bus.tvalid <= 1'b1;
                for (int b=0; b<egr_bus.DATA_BYTES; b++) begin
                    egr_bus.tdata[b*8 +: 8] <= send_data_buf[egr_port_rr][b*8 +: 8];
                end
                egr_bus.tuser  <= send_user_buf[egr_port_rr];
                dq_in_flight[egr_port_rr][0]                                             <= 1'b1;
                send_data_buf[egr_port_rr][0:MTU_BYTES*8-egr_bus.DATA_BYTES*8-1]         <= send_data_buf[egr_port_rr][egr_bus.DATA_BYTES*8:MTU_BYTES*8-1];
                send_data_buf[egr_port_rr][MTU_BYTES*8-egr_bus.DATA_BYTES*8:MTU_BYTES*8] <= '0;
                if (send_byte_length_buf[egr_port_rr] <= egr_bus.DATA_BYTES) begin
                    egr_bus.tlast                     <= 1'b1;
                    egr_bus.tkeep                     <= tkeep_comb;
                    send_byte_length_buf[egr_port_rr] <= 0;
                end else begin
                    send_byte_length_buf[egr_port_rr] <= send_byte_length_buf[egr_port_rr] - egr_bus.DATA_BYTES;
                end
            end
        end
    end


    ////////////////////////////////////////////////////////////////////////////////////////////////
    // SUB-SECTION:  Tx Packet Capture


    always_ff @(posedge core_clk_ifc.clk ) begin
        if (core_sreset_ifc.reset == core_sreset_ifc.ACTIVE_HIGH) begin
            tx_snoop_data_buf  <= '{default: '{default: '0}};
            tx_snoop_blen_buf  <= '{default: '{default: '0}};
            tx_snoop_wr_ptr    <= '{default: '0};
            send_packet_req_d  <= 1'b0;
        end else begin
            send_packet_req_d <= send_packet_req;
            if (send_packet_req && !send_packet_req_d) begin
                tx_snoop_data_buf[send_packet_user.egress_port][tx_snoop_wr_ptr[send_packet_user.egress_port]] <= send_packet_data;
                tx_snoop_blen_buf[send_packet_user.egress_port][tx_snoop_wr_ptr[send_packet_user.egress_port]] <= send_packet_byte_length;
                tx_snoop_wr_ptr[send_packet_user.egress_port]++;
            end
        end
    end


    ////////////////////////////////////////////////////////////////////////////////////////////////
    // SUB-SECTION: DUT


    p4_router_egress #(
        .NUM_8B_EGR_PHYS_PORTS  ( NUM_8B_PORTS      ),
        .NUM_16B_EGR_PHYS_PORTS ( NUM_16B_PORTS     ),
        .NUM_32B_EGR_PHYS_PORTS ( NUM_32B_PORTS     ),
        .NUM_64B_EGR_PHYS_PORTS ( NUM_64B_PORTS     ),
        .MTU_BYTES              ( MTU_BYTES         )
    ) DUT (
        .egr_bus                ( egr_bus               ),
        .egr_buf_ready          ( egr_buf_ready         ),
        .egr_8b_phys_ports      ( egr_8b_phys_ports     ),
        .egr_16b_phys_ports     ( egr_16b_phys_ports    ),
        .egr_32b_phys_ports     ( egr_32b_phys_ports    ),
        .egr_64b_phys_ports     ( egr_64b_phys_ports    ),
        .egr_phys_ports_enable  ( egr_phys_ports_enable ),
        .egr_cnts_clear         ( egr_cnts_clear        ),
        .egr_cnts               ( egr_cnts              ),
        .egr_ports_conneted     ( egr_ports_conneted    ),
        .egr_buf_full_drop      ( egr_buf_full_drop     )
    );

    // CDC

    `define DEF_CDC_FIFO(WIDTH)                                                         \
        axis_async_fifo_wrapper async_fifo (                                            \
            .axis_in             ( egr_``WIDTH``b_phys_ports[port_index]            ),  \
            .axis_out            ( egr_``WIDTH``b_phys_ports_cdc[port_index]        ),  \
            .axis_in_overflow    ( egr_``WIDTH``b_async_fifo_overflow[port_index]   ),  \
            .axis_in_bad_frame   (                                                  ),  \
            .axis_in_good_frame  (                                                  ),  \
            .axis_out_overflow   (                                                  ),  \
            .axis_out_bad_frame  (                                                  ),  \
            .axis_out_good_frame (                                                  )   \
        );

    generate
        for (genvar port_index=0; port_index<NUM_8B_PORTS; port_index++) begin : cdc_8b
            `DEF_CDC_FIFO(8);
        end
        for (genvar port_index=0; port_index<NUM_16B_PORTS; port_index++) begin : cdc_16b
            `DEF_CDC_FIFO(16);
        end
        for (genvar port_index=0; port_index<NUM_32B_PORTS; port_index++) begin : cdc_32b
            `DEF_CDC_FIFO(32);
        end
        for (genvar port_index=0; port_index<NUM_64B_PORTS; port_index++) begin : cdc_64b
            `DEF_CDC_FIFO(64);
        end
    endgenerate


    ////////////////////////////////////////////////////////////////////////////////////////////////
    // SUB-SECTION: Receive packet counter and demux verification


    // Modelsim didn't want to iterate over arrays of interfaces in an always_ff
    // pull tlast into a logic vector that Modelsim will allow iteration over.
    generate
        for (genvar i=0; i<NUM_8B_PORTS; i++) begin : axis_sigs_8b
            assign egr_phys_ports_tlast[EGR_PORT_INDEX_MAP[INDEX_8B][i]]  = egr_8b_phys_ports_cdc[i].tready & egr_8b_phys_ports_cdc[i].tvalid & egr_8b_phys_ports_cdc[i].tlast;
            assign egr_phys_ports_tvalid[EGR_PORT_INDEX_MAP[INDEX_8B][i]] = egr_8b_phys_ports_cdc[i].tready & egr_8b_phys_ports_cdc[i].tvalid & egr_8b_phys_ports_cdc[i].tvalid;
        end
        for (genvar i=0; i<NUM_16B_PORTS; i++) begin : axis_sigs_16b
            assign egr_phys_ports_tlast[EGR_PORT_INDEX_MAP[INDEX_16B][i]]  = egr_16b_phys_ports_cdc[i].tready & egr_16b_phys_ports_cdc[i].tvalid & egr_16b_phys_ports_cdc[i].tlast;
            assign egr_phys_ports_tvalid[EGR_PORT_INDEX_MAP[INDEX_16B][i]] = egr_16b_phys_ports_cdc[i].tready & egr_16b_phys_ports_cdc[i].tvalid & egr_16b_phys_ports_cdc[i].tvalid;
        end
        for (genvar i=0; i<NUM_32B_PORTS; i++) begin : axis_sigs_32b
            assign egr_phys_ports_tlast[EGR_PORT_INDEX_MAP[INDEX_32B][i]]  = egr_32b_phys_ports_cdc[i].tready & egr_32b_phys_ports_cdc[i].tvalid & egr_32b_phys_ports_cdc[i].tlast;
            assign egr_phys_ports_tvalid[EGR_PORT_INDEX_MAP[INDEX_32B][i]] = egr_32b_phys_ports_cdc[i].tready & egr_32b_phys_ports_cdc[i].tvalid & egr_32b_phys_ports_cdc[i].tvalid;
        end
        for (genvar i=0; i<NUM_64B_PORTS; i++) begin : axis_sigs_64b
            assign egr_phys_ports_tlast[EGR_PORT_INDEX_MAP[INDEX_64B][i]]  = egr_64b_phys_ports_cdc[i].tready & egr_64b_phys_ports_cdc[i].tvalid & egr_64b_phys_ports_cdc[i].tlast;
            assign egr_phys_ports_tvalid[EGR_PORT_INDEX_MAP[INDEX_64B][i]] = egr_64b_phys_ports_cdc[i].tready & egr_64b_phys_ports_cdc[i].tvalid & egr_64b_phys_ports_cdc[i].tvalid;
        end
    endgenerate

    always_ff @(posedge egr_port_clk_ifc.clk ) begin
        if (egr_port_sreset_ifc.reset == egr_port_sreset_ifc.ACTIVE_HIGH) begin
            received_count_array <= '{default: 0};
            received_count       <= 0;
            seq_cnt              <= 0;
            expected_egr_cnts    <= '{default: '{default: '{default: '0}}};
        end else begin
            packet_received <= 1'b0;
            for (int port=0; port<NUM_PORTS; port++) begin
                if (egr_phys_ports_tlast[port]) begin
                    if (verify_sequence) begin
                       `CHECK_EQUAL(port,seq_cnt % NUM_PORTS);
                        seq_cnt++;
                    end
                    received_count++;
                    packet_received <= 1'b1;
                    expected_egr_cnts[port][AXIS_PROFILE_PKT_CNT_INDEX]++;
                end
            end
        end
    end

    // Verify that there are no buffer overflows
    always_ff @( posedge core_clk_ifc.clk ) begin
        if (core_sreset_ifc.reset == core_sreset_ifc.ACTIVE_HIGH || egr_buf_full_drop_clear) begin
            egr_buf_full_drop_sticky <= '0;
        end else begin
            `CHECK_EQUAL(egr_buf_full_drop , 0);
            egr_buf_full_drop_sticky <= egr_buf_full_drop_sticky | egr_buf_full_drop;
        end
    end


    ////////////////////////////////////////////////////////////////////////////////////////////////
    // SUB-SECTION: Packet Sink and Check


    `define DEF_PKT_CHK(WIDTH)                                                                              \
        axis_array_packet_checker #(                                                                        \
            .NUM_PORTS                         ( NUM_``WIDTH``B_PORTS                                   ),  \
            .MODULE_ID_STRING_0                ( "Width Index"                                          ),  \
            .MODULE_ID_VALUE_0                 ( INDEX_``WIDTH``B                                       ),  \
            .MODULE_ID_STRING_1                ( "Array Index"                                          ),  \
            .AXIS_PACKET_IN_DATA_BYTES         ( egr_``WIDTH``b_phys_ports_cdc[0].DATA_BYTES            ),  \
            .AXIS_PACKET_IN_USER_WIDTH         ( egr_``WIDTH``b_phys_ports_cdc[0].USER_WIDTH            ),  \
            .AXIS_PACKET_IN_ALLOW_BACKPRESSURE ( egr_``WIDTH``b_phys_ports_cdc[0].ALLOW_BACKPRESSURE    ),  \
            .MTU_BYTES                         ( MTU_BYTES                                              ),  \
            .NUM_PACKETS_BEING_SENT            ( NUM_PACKETS_TO_SEND                                    )   \
        )  packet_checker_``WIDTH``b  (                                                                     \
            .axis_packet_in ( egr_``WIDTH``b_phys_ports_cdc                                     ),          \
            .num_tx_pkts    ( tx_snoop_wr_ptr[EGR_``WIDTH``B_START +: NUM_``WIDTH``B_PORTS]     ),          \
            .expected_pkts  ( tx_snoop_data_buf[EGR_``WIDTH``B_START +: NUM_``WIDTH``B_PORTS]   ),          \
            .expected_blens ( tx_snoop_blen_buf[EGR_``WIDTH``B_START +: NUM_``WIDTH``B_PORTS]   ),          \
            .expected_dests ( '{default: '{default: '0}}                                        )           \
        );

    generate
        if (NUM_8B_PORTS) begin : packet_checker_8b_g
            `DEF_PKT_CHK(8);
        end

        if (NUM_16B_PORTS) begin : packet_checker_16b_g
            `DEF_PKT_CHK(16);
        end

        if (NUM_32B_PORTS) begin : packet_checker_32b_g
            `DEF_PKT_CHK(32);
        end

        if (NUM_64B_PORTS) begin : packet_checker_64b_g
            `DEF_PKT_CHK(64);
        end
    endgenerate


    ////////////////////////////////////////////////////////////////////////////////////////////////
    // SUB-SECTION: Verify that there are no buffer overflows


    always_ff @( posedge core_clk_ifc.clk ) begin
        if (core_sreset_ifc.reset != core_sreset_ifc.ACTIVE_HIGH) begin
            `CHECK_EQUAL(egr_8b_async_fifo_overflow , 0);
            `CHECK_EQUAL(egr_16b_async_fifo_overflow , 0);
            `CHECK_EQUAL(egr_32b_async_fifo_overflow , 0);
            `CHECK_EQUAL(egr_64b_async_fifo_overflow , 0);
        end
    end


    ////////////////////////////////////////////////////////////////////////////////////////////////
    // SECTION: Tasks


    task automatic send_packet (
        input int                     send_packet_port,
        input bit [MTU_BYTES_LOG-1:0] packet_byte_length
    ); begin
            // Wait till we can send data
            @(posedge core_clk_ifc.clk && !send_packet_busy[send_packet_port]);
            #1;
            send_packet_user.egress_port = send_packet_port;
            send_packet_byte_length      = packet_byte_length;
            axis_packet_formatter #( EGR_AXIS_DATA_BYTES,  MAX_PKT_EGR_WLEN , MTU_BYTES)::get_packet(PAYLOAD_TYPE, packet_byte_length, send_packet_data);
            send_packet_req = 1'b1;
            @(posedge core_clk_ifc.clk);
            #1;
            send_packet_req = 1'b0;
        end
    endtask;

    task automatic send_random_length_packet (
        input int send_packet_port
    ); begin
            send_packet(send_packet_port, $urandom_range(PACKET_MAX_BLEN, PACKET_MIN_BLEN));
       end
    endtask

    task automatic check_packet_counts();
        begin
            // Compare tx and rx counts
            `CHECK_EQUAL(received_count, expected_count);
            for (int i=0; i<NUM_PORTS; i++) begin
                // Check that the expected number of packets were counted by the DUT egress counters
                `CHECK_EQUAL(egr_cnts[i][AXIS_PROFILE_PKT_CNT_INDEX], expected_egr_cnts[i][AXIS_PROFILE_PKT_CNT_INDEX]);
                // Verify that the DUT egress counters clears and don't disrupt other counts
                egr_cnts_clear[i] = 1'b1;
                @(posedge core_clk_ifc.clk);
                #1;
                `CHECK_EQUAL(egr_cnts[i][AXIS_PROFILE_PKT_CNT_INDEX], 0);
            end
        end
    endtask


    ////////////////////////////////////////////////////////////////////////////////////////////////
    // SECTION: Tests


    `TEST_SUITE begin
        `TEST_SUITE_SETUP begin
            $timeformat(-9, 3, " ns", 20);
            core_clk_ifc.clk     = 1'b0;
            egr_port_clk_ifc.clk = 1'b0;
            send_packet_req      = 1'b0;
        end

        `TEST_CASE_SETUP begin
            egr_cnts_clear = '1;
            @(posedge core_clk_ifc.clk);
            #1;
            egr_cnts_clear = '0;

            egr_phys_ports_enable   = '1;
            egr_buf_full_drop_clear = 1'b0;
            send_packet_req         = 1'b0;
            verify_sequence         = 1'b0;
            expected_count          = NUM_PACKETS_TO_SEND;

            core_sreset_ifc.reset     = core_sreset_ifc.ACTIVE_HIGH;
            egr_port_sreset_ifc.reset = egr_port_sreset_ifc.ACTIVE_HIGH;

            repeat (10) @(posedge egr_port_clk_ifc.clk);
            egr_port_sreset_ifc.reset = ~egr_port_sreset_ifc.ACTIVE_HIGH;
            @(posedge core_clk_ifc.clk);
            core_sreset_ifc.reset = ~core_sreset_ifc.ACTIVE_HIGH;
            repeat (8) @(posedge core_clk_ifc.clk);
        end

        // Send packets to all ports
        `TEST_CASE("send_to_all_ports") begin

            automatic bit egress_active = 1'b1;

            expected_count = NUM_PACKETS_TO_SEND;

            for (int pkt=0; pkt<NUM_PACKETS_TO_SEND; pkt++) begin
                // Send random length packet to each port sequentially
                send_random_length_packet(pkt % NUM_PORTS);
            end

            // wait for packets to exit the DUT
            while (egress_active) begin
                egress_active = 1'b0;
                for (int i=0; i<64; i++) begin
                    @(posedge egr_port_clk_ifc.clk);
                    #1;
                    egress_active = egress_active | |egr_phys_ports_tvalid;
                end
            end
            repeat (MAX_PKT_WLEN_8B) @(posedge egr_port_clk_ifc.clk);
            @(core_clk_ifc.clk);

            check_packet_counts;
        end

        // Send packets with all ports disabled
        `TEST_CASE("disable_all_ports") begin
            automatic bit egress_active = 1'b1;

            egr_phys_ports_enable = '0;
            expected_count = 0;

            for (int pkt=0; pkt<NUM_PACKETS_TO_SEND; pkt++) begin
                send_random_length_packet(pkt % NUM_PORTS);
            end

            // wait for packets to exit the DUT
            while (egress_active) begin
                egress_active = 1'b0;
                for (int i=0; i<64; i++) begin
                    @(posedge egr_port_clk_ifc.clk);
                    #1;
                    egress_active = egress_active | |egr_phys_ports_tvalid;
                end
            end

            check_packet_counts;
        end

        // Send packets with one port disabled
        `TEST_CASE("disable_one_port") begin
            automatic int disabled_port = $urandom() % NUM_PORTS;
            automatic int port;
            automatic bit egress_active = 1'b1;

            egr_phys_ports_enable[disabled_port] = 1'b0;
            expected_count = 0;

            for (int pkt=0; pkt<NUM_PACKETS_TO_SEND; pkt++) begin
                port = pkt % NUM_PORTS;
                if (port != disabled_port) expected_count += 1;
                send_random_length_packet(pkt % NUM_PORTS);
            end

            // wait for packets to exit the DUT
            while (egress_active) begin
                egress_active = 1'b0;
                for (int i=0; i<64; i++) begin
                    @(posedge egr_port_clk_ifc.clk);
                    #1;
                    egress_active = egress_active | |egr_phys_ports_tvalid;
                end
            end

            check_packet_counts;
        end
    end

    `WATCHDOG(10ms);

endmodule
