// CONFIDENTIAL
// Copyright (c) 2024 Kepler Communications Inc.

/**
 * MPLS Router Package
**/

package mpls_router_pkg;



endpackage