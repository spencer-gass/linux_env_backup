// CONFIDENTIAL
// Copyright (c) 2024 Kepler Communications Inc.

/**
 * P4 Router Package
**/

`default_nettype none

package p4_router_pkg;

    ////////////////////////////////////////////////////////////////////////////////////////////////
    // SECTION: ENUMs

    enum {
        RESERVED,
        ECHO_PHYS_PORT,
        FRR_T1_ECP,
        NUM_VNP4_IP_OPTIONS
    } vnp4_ip_options;

    enum {
        INDEX_8B,
        INDEX_16B,
        INDEX_32B,
        INDEX_64B,
        NUM_AXIS_ARRAYS
    } port_width_indecies;

    enum {
        GREEN,
        YELLOW,
        RED,
        UNCOLORED,
        NUM_POLICER_COLORS
    } policer_colors;


    ////////////////////////////////////////////////////////////////////////////////////////////////
    // SECTION: Physical Port Array Related Constants and Functions

    localparam int NUM_ING_AXIS_ARRAYS = NUM_AXIS_ARRAYS;
    localparam int NUM_EGR_AXIS_ARRAYS = NUM_AXIS_ARRAYS;

    function int get_max_num_ports_per_array(
        input int array [NUM_AXIS_ARRAYS-1:0]
    );
        automatic int max = 0;
        for (int i=0; i<NUM_AXIS_ARRAYS; i++) begin
            if (array[i] > max) begin
                max = array[i];
            end
        end
        return max;
    endfunction


    ////////////////////////////////////////////////////////////////////////////////////////////////
    // SECTION: Stats Counters

    localparam int AXIS_PROFILE_BYTE_CNT_INDEX  = 0;
    localparam int AXIS_PROFILE_PKT_CNT_INDEX   = 5;
    localparam int AXIS_PROFILE_ERR_CNT_INDEX   = 6;

    localparam int ING_COUNTERS_WIDTH = 32;
    localparam int EGR_COUNTERS_WIDTH = 32;


    ////////////////////////////////////////////////////////////////////////////////////////////////
    // SECTION: Metadata structs Conveyed By AXIS.tuser

    localparam INGRESS_METADATA_INGRESS_PORT_WIDTH = 5;
    localparam VNP4_WRAPPER_METADATA_EGRESS_PORT_WIDTH = 5;

    typedef struct packed {
        logic [INGRESS_METADATA_INGRESS_PORT_WIDTH-1:0]  ingress_port;
    } ingress_metadata_t;

    typedef struct packed {
        logic [INGRESS_METADATA_INGRESS_PORT_WIDTH-1:0]  ingress_port;
        logic [VNP4_WRAPPER_METADATA_EGRESS_PORT_WIDTH-1:0]  egress_port;
        logic [2:0]  prio;
        logic [13:0] byte_length;
    } vnp4_wrapper_metadata_t;

    typedef struct packed {
        logic [INGRESS_METADATA_INGRESS_PORT_WIDTH-1:0]  ingress_port;
        logic [VNP4_WRAPPER_METADATA_EGRESS_PORT_WIDTH-1:0]  egress_port;
        logic [2:0]  prio;
        logic [13:0] byte_length;
        logic [1:0]  policer_color;
    } policer_metadata_t;

    typedef struct packed {
        logic [15:0]  tail_ptr;
        logic [15:0]  current_page_ptr;
        logic [15:0]  next_page_ptr;
    } cong_man_metadata_t;

    typedef struct packed {
        logic [VNP4_WRAPPER_METADATA_EGRESS_PORT_WIDTH-1:0]  egress_port;
    } queue_system_metadata_t;

    localparam int INGRESS_METADATA_WIDTH = $bits(ingress_metadata_t);
    localparam int VNP4_WRAPPER_METADATA_WIDTH = $bits(vnp4_wrapper_metadata_t);
    localparam int POLICER_METADATA_WIDTH = $bits(policer_metadata_t);
    localparam int CONG_MAN_METADATA_WIDTH = $bits(cong_man_metadata_t);
    localparam int QUEUE_SYS_METADATA_WIDTH = $bits(queue_system_metadata_t);


    ////////////////////////////////////////////////////////////////////////////////////////////////
    // SECTION: Queue System

    localparam int POLICER_COLOR_BITS = 2;
    localparam int PRIO_BITS = 3;

    function policer_metadata_t add_policer_color_to_metadata(
        input logic [POLICER_COLOR_BITS-1:0] policer_color,
        input vnp4_wrapper_metadata_t vnp4_wrapper_metadata
    );
        automatic policer_metadata_t policer_metadata;

        policer_metadata.ingress_port = vnp4_wrapper_metadata.ingress_port;
        policer_metadata.egress_port  = vnp4_wrapper_metadata.egress_port;
        policer_metadata.prio         = vnp4_wrapper_metadata.prio;
        policer_metadata.byte_length  = vnp4_wrapper_metadata.byte_length;
        policer_metadata.policer_color = policer_color;

        return policer_metadata;
    endfunction

    localparam int NUM_QUEUES_PER_EGR_PORT = 4;
    localparam int NUM_QUEUES_PER_EGR_PORT_LOG = $clog2(NUM_QUEUES_PER_EGR_PORT);
    localparam int DQ_LATENCY = 4; // cycles between scheduler dequeue request and dequeue notification
    localparam int POLICER_TABLE_WIDTH = 64; /// revisit when you design the policer
    localparam int DROP_THRESH_TABLE_WIDTH = 3*22; // 3xMAX_QUEUE_OCCUPANCY_LOG


    ////////////////////////////////////////////////////////////////////////////////////////////////
    // SECTION: Metadata Structs Conveyed Over AXI4Lite.rdata and AXI4Lite.wdata

    // Used for AXI4Lite rdata and wdata, so keep total bit-width byte-alligned.
    typedef struct packed {
        logic [15:0] tail_ptr;
        logic [14:0] current_page_ptr;
        logic        current_page_valid;
    } queue_tail_pointer_read_t;

    typedef struct packed {
        logic [15:0] new_tail_ptr;
        logic [14:0] next_page_ptr;
        logic        malloc_approved;
    } queue_tail_pointer_write_t;

    localparam QUEUE_TAIL_POINTER_DATALEN = 32;

    typedef struct packed {
        logic [15:0] head_ptr;
        logic [15:0] page_ptr;
    } queue_head_pointer_read_t;

    localparam QUEUE_HEAD_POINTER_DATALEN = 32;


endpackage

`default_nettype wire